library ieee;
use ieee.std_logic_1164.all;

entity pipes is
	generic(
		--Nisam siguran da li sam dobro izracunao opseg
		C_LAST_POS : integer := (2*(1023 - 72) + 64 + 72);
		
		C_FIRST_POS : integer range 1023 to C_LAST_POS; 	-- Initial position of a pipe.
		C_NEXT_POS 	: integer range 1023 to C_LAST_POS;		-- Position on wich pipe goes after reaching left border of a display.
		
		C_PIPE_WIDTH	: integer := 64;
		C_WINDOW_WIDTH	: integer := 32;
		
		C_PIPE_VELOCITY	: integer := 1;
		
		H_DISPLAY	: integer := 1024;
		V_DISPLAY	: integer := 768
	);
	port(
		clk65M				: in std_logic;							-- clock 65Mhz
		reset				: in std_logic; 						-- reset
		started				: in std_logic;							-- if game is on or off
		hpos 				: in integer range 0 to H_DISPLAY - 1;	-- output of vga_controller
		vpos 				: in integer range 0 to V_DISPLAY - 1;	-- output of vga_controller
		ref_tick			: in std_logic;							-- output of vga_controller
		window_ypos			: in integer range 32 to 735;			-- y position of a window
		--pipe_xpos			: out integer range -C_PIPE_WIDTH to (C_LAST_POS + C_PIPE_WIDTH);
		Rout, Gout, Bout	: out std_logic_vector(7 downto 0)		-- input in vga_controller
	);
end pipes;

architecture Behavioral of pipes is

	constant BCKG_COLOR : std_logic_vector(23 downto 0) := x"777777";
	constant PIPE_COLOR : std_logic_vector(23 downto 0) := x"007700";

	signal xpos		: integer range -C_PIPE_WIDTH to (C_LAST_POS + C_PIPE_WIDTH);
	signal on_pipe	: std_logic;
	signal color 	: std_logic_vector(23 downto 0);

begin
	
	-- Update position. If reset is active or game is
	-- not on then the position of the pipe has initial value. 
	-- Otherwise on rising clock edge on the end of the frame if pipe
	-- reached right edge of the display the position of the pipe is set
	-- to be on right edge of the display. If pipe did not reached left edge,
	-- position of the pipe is decremented by defined constant.
	process(clk65M, reset, ref_tick, started) is
	begin
		if reset = '1' or started = '0' then
			xpos <= C_FIRST_POS;
		else
			if rising_edge(clk65M) then
				if ref_tick = '1' then
					if xpos < -C_PIPE_WIDTH then
						xpos <= C_NEXT_POS;
					else  
						xpos <= xpos - C_PIPE_VELOCITY;
					end if;
				end if;
			end if;
		end if;
	end process;
	
	--pipe_xpos <= xpos;
	
	-- If vpos and hpos are on the pipe, signal on_pipe is active.
	on_pipe <= '1' when ((hpos >= xpos and hpos < (xpos + C_PIPE_WIDTH)) and (vpos <= window_ypos and vpos > (window_ypos + C_WINDOW_WIDTH))) else
					'0';
	
	-- If reset is active color of every pixel is black.
	-- If signal on_pipe is active, color that goes to the vga_controller 
	-- is the color of the pipe. If not, color is color of background.
	process(reset, on_pipe) is
	begin
		if reset = '1' then 
			color <= (others => '0');
		else
			if on_pipe = '1' then
				color <= PIPE_COLOR;
			else
				color <= BCKG_COLOR;
			end if;
		end if;
	end process;
	
	Rout <= color(23 downto 16);
	Gout <= color(15 downto 8);
	Bout <= color(7 downto 0);

end Behavioral;